-- George Landis
-- Lab 02
-- ECET 109

library ieee; -- allows the use of all ieee libraries
use ieee.std_logic_1164.all; -- contains definitions of types, subtypes and functions
use ieee.numeric_std.all; -- numeric types and arthmetic functions for use with synthesis tools

entity Lab_02 is
-- in this area you will define the inputs and outputs for the circuit.

end entity;

architecture learning_VHDL of Lab_02 is -- the text "learning_VHDL" can be any name you like
begin -- all architecture statements use the key word begin to identify the starting point of the logic

end learning_VHDL;-- all architecture statements use the key word "end" to denote the stoping point.


